library ieee;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use STD.TEXTIO.ALL;

entity mem_instruct is
    port(
        PC: in std_logic_vector(31 downto 0);-- entree d'adresse
        instr: out std_logic_vector(31 downto 0)
    );
end mem_instruct;

architecture behavioral of mem_instruct is
    -- Declaration du tableau memoire
    type mem_array is array(0 to 63) of std_logic_vector(31 downto 0);
    signal mem : mem_array := ("11100000010000000000000000000000", 
                               "11100010100000000010000000000101", 
                               "11100010100000000011000000001100",
                               "11100010010000110111000000001001",
                               "11100001100001110100000000000010",
                               "11100000000000110101000000000100",
                               "11100000100001010101000000000100",
                               "11100000010101011000000000000111",
                               "11100000010100111000000000000100",
                               "11100010100000000101000000000000",
                               "11100000010101111000000000000010",
                               "10110010100001010111000000000001",
                               "11100000010001110111000000000010",
                               "11100101100000110111000001010100",
                               "11100101100100000010000001100000",
                               "11100000100010000101000000000000",
                               "11100010100000000010000000001110",
                               "11100010100000000010000000001101",
                               "11100010100000000010000000001010",
                               "11100101100000000010000001100100",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               -- 32 �l�ments suppl�mentaires pour compl�ter le tableau (indices 32 � 63)
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000",
                               "00000000000000000000000000000000");
begin
    -- Lecture en tout temps
    instr <= mem(TO_INTEGER(unsigned(PC(6 downto 2))));
    
end behavioral;